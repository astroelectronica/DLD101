.title KiCad schematic
.include "C:/AE/DLD101/_models/2N7002.spice.txt"
.include "C:/AE/DLD101/_models/DLD101.spice.txt"
.include "C:/AE/DLD101/_models/XPE_SPICE.lib"
R3 VCC /D {RD}
R2 /G 0 {RPD}
R1 /DIM /G {RG}
V1 /DIM 0 PULSE(0 {VPUL} {DELAY} {TR} {TF} {DUTY} {CYCLE})
D4 /L3 /L4 XLampXPEblue
D3 /L2 /L3 XLampXPEblue
D2 /L1 /L2 XLampXPEblue
D1 VCC /L1 XLampXPEblue
R4 /SET 0 {RSET}
XU2 /K /D /D 0 unconnected-_U2-R1-PadP6_ /SET /SET DLD101
D7 /L6 /L7 XLampXPEblue
D8 /L7 /K XLampXPEblue
D6 /L5 /L6 XLampXPEblue
D5 /L4 /L5 XLampXPEblue
XQ1 /D /G 0 N7002
V2 VCC 0 {VSOURCE}
.end
