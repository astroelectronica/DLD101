.title KiCad schematic
.include "C:/AE/DLD101/_models/2N7002.spice.txt"
.include "C:/AE/DLD101/_models/DLD101.spice.txt"
.include "C:/AE/DLD101/_models/XPE_SPICE.lib"
R3 VCC /D {RD}
R2 /G 0 {RPD}
R1 /DIM /G {RG}
V1 /DIM 0 PULSE(0 {VPUL} {DELAY} {TR} {TF} {DUTY} {CYCLE})
D4 /L3 /L4 XLampXPEgreen
D3 /L2 /L3 XLampXPEgreen
D2 /L1 /L2 XLampXPEgreen
D1 VCC /L1 XLampXPEgreen
R4 /SET 0 {RSET}
XU2 /K /D /D 0 unconnected-_U2-R1-PadP6_ /SET /SET DLD101
D7 /L6 /L7 XLampXPEgreen
D8 /L7 /K XLampXPEgreen
D6 /L5 /L6 XLampXPEgreen
D5 /L4 /L5 XLampXPEgreen
XQ1 /D /G 0 N7002
V2 VCC 0 {VSOURCE}
.end
